magic
tech sky130A
magscale 1 2
timestamp 1713492000
<< poly >>
rect 17293 7100 18108 7202
rect 18006 6660 18108 7100
rect 17910 6640 18125 6660
rect 17910 6509 17930 6640
rect 18100 6509 18125 6640
rect 17910 6490 18125 6509
<< polycont >>
rect 17930 6509 18100 6640
<< locali >>
rect 17910 6640 18125 6660
rect 17910 6509 17930 6640
rect 18100 6509 18125 6640
rect 17910 6490 18125 6509
rect 18468 6253 18801 6660
rect 19169 6541 19430 6647
rect 18468 6120 18523 6253
rect 18736 6120 18801 6253
rect 18468 6086 18801 6120
<< viali >>
rect 17930 6509 18100 6640
rect 18523 6120 18736 6253
<< metal1 >>
rect 17910 6640 18125 6660
rect 17910 6509 17930 6640
rect 18100 6509 18125 6640
rect 17910 6490 18125 6509
rect 18468 6253 18801 6298
rect 18468 6120 18523 6253
rect 18736 6120 18801 6253
rect 18468 6086 18801 6120
<< via1 >>
rect 17930 6509 18100 6640
rect 18523 6120 18736 6253
<< metal2 >>
rect 17910 6640 18125 6660
rect 17910 6509 17930 6640
rect 18100 6509 18125 6640
rect 17910 6490 18125 6509
rect 18468 6253 18801 6298
rect 18468 6120 18523 6253
rect 18736 6120 18801 6253
rect 18468 6086 18801 6120
<< via2 >>
rect 17930 6509 18100 6640
rect 18523 6120 18736 6253
rect 16026 3693 16303 3959
rect 23658 3672 23828 3838
<< metal3 >>
rect 17910 6640 18125 6660
rect 17910 6509 17930 6640
rect 18100 6509 18125 6640
rect 17910 6490 18125 6509
rect 18468 6253 18801 6298
rect 18468 6120 18523 6253
rect 18736 6120 18801 6253
rect 18468 6086 18801 6120
rect 17200 4672 17449 5155
rect 17200 4500 17224 4672
rect 17418 4500 17449 4672
rect 17200 4451 17449 4500
rect 15967 3959 16366 4023
rect 15967 3693 16026 3959
rect 16303 3693 16366 3959
rect 15967 3619 16366 3693
rect 23544 3838 23944 3864
rect 23544 3672 23658 3838
rect 23828 3672 23944 3838
rect 23544 3606 23944 3672
<< via3 >>
rect 20640 7687 20788 7827
rect 17930 6509 18100 6640
rect 18523 6120 18736 6253
rect 17224 4500 17418 4672
rect 16026 3693 16303 3959
rect 23658 3672 23828 3838
<< metal4 >>
rect 798 44952 858 45152
rect 1534 44952 1594 45152
rect 2270 44952 2330 45152
rect 3006 44952 3066 45152
rect 3742 44952 3802 45152
rect 4478 44952 4538 45152
rect 5214 44952 5274 45152
rect 5950 44952 6010 45152
rect 6686 44952 6746 45152
rect 7422 44952 7482 45152
rect 8158 44952 8218 45152
rect 8894 44952 8954 45152
rect 9630 44952 9690 45152
rect 10366 44952 10426 45152
rect 11102 44952 11162 45152
rect 11838 44952 11898 45152
rect 12574 44952 12634 45152
rect 13310 44952 13370 45152
rect 14046 44952 14106 45152
rect 14782 44952 14842 45152
rect 15518 44952 15578 45152
rect 16254 44952 16314 45152
rect 16990 44952 17050 45152
rect 17726 44952 17786 45152
rect 18462 44952 18522 45152
rect 19198 44952 19258 45152
rect 19934 44952 19994 45152
rect 20670 44952 20730 45152
rect 21406 44952 21466 45152
rect 22142 44952 22202 45152
rect 22878 44952 22938 45152
rect 23614 44952 23674 45152
rect 24350 44952 24410 45152
rect 25086 44952 25146 45152
rect 25822 44952 25882 45152
rect 26558 44952 26618 45152
rect 27294 44952 27354 45152
rect 28030 44952 28090 45152
rect 28766 44952 28826 45152
rect 29502 44952 29562 45152
rect 30238 44952 30298 45152
rect 30974 44952 31034 45152
rect 31710 44952 31770 45152
rect 200 1000 500 44152
rect 9800 6803 10100 44152
rect 20599 7827 20822 7877
rect 20599 7687 20640 7827
rect 20788 7687 20822 7827
rect 9635 6022 16926 6803
rect 17910 6640 18125 6660
rect 17910 6509 17930 6640
rect 18100 6509 18125 6640
rect 9800 1000 10100 6022
rect 17910 5849 18125 6509
rect 18468 6253 19430 6290
rect 18468 6120 18523 6253
rect 18736 6120 19430 6253
rect 18468 6086 19430 6120
rect 17910 5621 18549 5849
rect 17185 4672 17476 4726
rect 17185 4500 17224 4672
rect 17418 4500 17476 4672
rect 17185 4068 17476 4500
rect 11977 3959 16385 4022
rect 11977 3693 16026 3959
rect 16303 3693 16385 3959
rect 11977 3618 16385 3693
rect 12078 435 12281 3618
rect 17222 1348 17438 4068
rect 18262 3121 18546 5621
rect 18018 2908 18546 3121
rect 13600 1132 17438 1348
rect 9232 315 12281 435
rect 400 0 520 200
rect 4816 0 4936 200
rect 9232 0 9352 315
rect 12078 274 12281 315
rect 13648 0 13768 1132
rect 18064 0 18184 2908
rect 18262 2872 18546 2908
rect 19169 1930 19429 6086
rect 20599 2790 20822 7687
rect 23544 3862 23942 3864
rect 23544 3838 31494 3862
rect 23544 3672 23658 3838
rect 23828 3672 31494 3838
rect 23544 3618 31494 3672
rect 23544 3606 23942 3618
rect 20599 2567 27068 2790
rect 19169 1716 22647 1930
rect 19169 1693 19429 1716
rect 22480 0 22600 1716
rect 26896 0 27016 2567
rect 31312 0 31432 3618
use opamp  opamp_0 ~/Desktop/opamp/layout
timestamp 1713491752
transform 1 0 21146 0 1 8051
box -5777 -4445 2796 16960
<< labels >>
flabel metal4 s 30974 44952 31034 45152 0 FreeSans 480 90 0 0 clk
port 0 nsew signal input
flabel metal4 s 31710 44952 31770 45152 0 FreeSans 480 90 0 0 ena
port 1 nsew signal input
flabel metal4 s 30238 44952 30298 45152 0 FreeSans 480 90 0 0 rst_n
port 2 nsew signal input
flabel metal4 s 31312 0 31432 200 0 FreeSans 960 0 0 0 ua[0]
port 3 nsew signal bidirectional
flabel metal4 s 26896 0 27016 200 0 FreeSans 960 0 0 0 ua[1]
port 4 nsew signal bidirectional
flabel metal4 s 22480 0 22600 200 0 FreeSans 960 0 0 0 ua[2]
port 5 nsew signal bidirectional
flabel metal4 s 18064 0 18184 200 0 FreeSans 960 0 0 0 ua[3]
port 6 nsew signal bidirectional
flabel metal4 s 13648 0 13768 200 0 FreeSans 960 0 0 0 ua[4]
port 7 nsew signal bidirectional
flabel metal4 s 9232 0 9352 200 0 FreeSans 960 0 0 0 ua[5]
port 8 nsew signal bidirectional
flabel metal4 s 4816 0 4936 200 0 FreeSans 960 0 0 0 ua[6]
port 9 nsew signal bidirectional
flabel metal4 s 400 0 520 200 0 FreeSans 960 0 0 0 ua[7]
port 10 nsew signal bidirectional
flabel metal4 s 29502 44952 29562 45152 0 FreeSans 480 90 0 0 ui_in[0]
port 11 nsew signal input
flabel metal4 s 28766 44952 28826 45152 0 FreeSans 480 90 0 0 ui_in[1]
port 12 nsew signal input
flabel metal4 s 28030 44952 28090 45152 0 FreeSans 480 90 0 0 ui_in[2]
port 13 nsew signal input
flabel metal4 s 27294 44952 27354 45152 0 FreeSans 480 90 0 0 ui_in[3]
port 14 nsew signal input
flabel metal4 s 26558 44952 26618 45152 0 FreeSans 480 90 0 0 ui_in[4]
port 15 nsew signal input
flabel metal4 s 25822 44952 25882 45152 0 FreeSans 480 90 0 0 ui_in[5]
port 16 nsew signal input
flabel metal4 s 25086 44952 25146 45152 0 FreeSans 480 90 0 0 ui_in[6]
port 17 nsew signal input
flabel metal4 s 24350 44952 24410 45152 0 FreeSans 480 90 0 0 ui_in[7]
port 18 nsew signal input
flabel metal4 s 23614 44952 23674 45152 0 FreeSans 480 90 0 0 uio_in[0]
port 19 nsew signal input
flabel metal4 s 22878 44952 22938 45152 0 FreeSans 480 90 0 0 uio_in[1]
port 20 nsew signal input
flabel metal4 s 22142 44952 22202 45152 0 FreeSans 480 90 0 0 uio_in[2]
port 21 nsew signal input
flabel metal4 s 21406 44952 21466 45152 0 FreeSans 480 90 0 0 uio_in[3]
port 22 nsew signal input
flabel metal4 s 20670 44952 20730 45152 0 FreeSans 480 90 0 0 uio_in[4]
port 23 nsew signal input
flabel metal4 s 19934 44952 19994 45152 0 FreeSans 480 90 0 0 uio_in[5]
port 24 nsew signal input
flabel metal4 s 19198 44952 19258 45152 0 FreeSans 480 90 0 0 uio_in[6]
port 25 nsew signal input
flabel metal4 s 18462 44952 18522 45152 0 FreeSans 480 90 0 0 uio_in[7]
port 26 nsew signal input
flabel metal4 s 5950 44952 6010 45152 0 FreeSans 480 90 0 0 uio_oe[0]
port 27 nsew signal output
flabel metal4 s 5214 44952 5274 45152 0 FreeSans 480 90 0 0 uio_oe[1]
port 28 nsew signal output
flabel metal4 s 4478 44952 4538 45152 0 FreeSans 480 90 0 0 uio_oe[2]
port 29 nsew signal output
flabel metal4 s 3742 44952 3802 45152 0 FreeSans 480 90 0 0 uio_oe[3]
port 30 nsew signal output
flabel metal4 s 3006 44952 3066 45152 0 FreeSans 480 90 0 0 uio_oe[4]
port 31 nsew signal output
flabel metal4 s 2270 44952 2330 45152 0 FreeSans 480 90 0 0 uio_oe[5]
port 32 nsew signal output
flabel metal4 s 1534 44952 1594 45152 0 FreeSans 480 90 0 0 uio_oe[6]
port 33 nsew signal output
flabel metal4 s 798 44952 858 45152 0 FreeSans 480 90 0 0 uio_oe[7]
port 34 nsew signal output
flabel metal4 s 11838 44952 11898 45152 0 FreeSans 480 90 0 0 uio_out[0]
port 35 nsew signal output
flabel metal4 s 11102 44952 11162 45152 0 FreeSans 480 90 0 0 uio_out[1]
port 36 nsew signal output
flabel metal4 s 10366 44952 10426 45152 0 FreeSans 480 90 0 0 uio_out[2]
port 37 nsew signal output
flabel metal4 s 9630 44952 9690 45152 0 FreeSans 480 90 0 0 uio_out[3]
port 38 nsew signal output
flabel metal4 s 8894 44952 8954 45152 0 FreeSans 480 90 0 0 uio_out[4]
port 39 nsew signal output
flabel metal4 s 8158 44952 8218 45152 0 FreeSans 480 90 0 0 uio_out[5]
port 40 nsew signal output
flabel metal4 s 7422 44952 7482 45152 0 FreeSans 480 90 0 0 uio_out[6]
port 41 nsew signal output
flabel metal4 s 6686 44952 6746 45152 0 FreeSans 480 90 0 0 uio_out[7]
port 42 nsew signal output
flabel metal4 s 17726 44952 17786 45152 0 FreeSans 480 90 0 0 uo_out[0]
port 43 nsew signal output
flabel metal4 s 16990 44952 17050 45152 0 FreeSans 480 90 0 0 uo_out[1]
port 44 nsew signal output
flabel metal4 s 16254 44952 16314 45152 0 FreeSans 480 90 0 0 uo_out[2]
port 45 nsew signal output
flabel metal4 s 15518 44952 15578 45152 0 FreeSans 480 90 0 0 uo_out[3]
port 46 nsew signal output
flabel metal4 s 14782 44952 14842 45152 0 FreeSans 480 90 0 0 uo_out[4]
port 47 nsew signal output
flabel metal4 s 14046 44952 14106 45152 0 FreeSans 480 90 0 0 uo_out[5]
port 48 nsew signal output
flabel metal4 s 13310 44952 13370 45152 0 FreeSans 480 90 0 0 uo_out[6]
port 49 nsew signal output
flabel metal4 s 12574 44952 12634 45152 0 FreeSans 480 90 0 0 uo_out[7]
port 50 nsew signal output
flabel metal4 200 1000 500 44152 1 FreeSans 2 0 0 0 VPWR
port 51 nsew power bidirectional
flabel metal4 9800 1000 10100 44152 1 FreeSans 2 0 0 0 VGND
port 52 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 32200 45152
<< end >>
