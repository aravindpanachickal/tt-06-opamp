VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO tt_um_duk_opamp
  CLASS BLOCK ;
  FOREIGN tt_um_duk_opamp ;
  ORIGIN 0.000 0.000 ;
  SIZE 161.000 BY 225.760 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 154.870 224.760 155.170 225.760 ;
    END
  END clk
  PIN ena
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 158.550 224.760 158.850 225.760 ;
    END
  END ena
  PIN rst_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 151.190 224.760 151.490 225.760 ;
    END
  END rst_n
  PIN ua[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 28.808649 ;
    PORT
      LAYER met4 ;
        RECT 156.560 0.000 157.160 1.000 ;
    END
  END ua[0]
  PIN ua[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 8.410000 ;
    PORT
      LAYER met4 ;
        RECT 134.480 0.000 135.080 1.000 ;
    END
  END ua[1]
  PIN ua[2]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 28.500000 ;
    PORT
      LAYER met4 ;
        RECT 112.400 0.000 113.000 1.000 ;
    END
  END ua[2]
  PIN ua[3]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 28.500000 ;
    PORT
      LAYER met4 ;
        RECT 90.320 0.000 90.920 1.000 ;
    END
  END ua[3]
  PIN ua[4]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.215000 ;
    PORT
      LAYER met4 ;
        RECT 68.240 0.000 68.840 1.000 ;
    END
  END ua[4]
  PIN ua[5]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.700000 ;
    ANTENNADIFFAREA 289.766205 ;
    PORT
      LAYER met4 ;
        RECT 46.160 0.000 46.760 1.000 ;
    END
  END ua[5]
  PIN ua[6]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 24.080 0.000 24.680 1.000 ;
    END
  END ua[6]
  PIN ua[7]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 2.000 0.000 2.600 1.000 ;
    END
  END ua[7]
  PIN ui_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 147.510 224.760 147.810 225.760 ;
    END
  END ui_in[0]
  PIN ui_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 143.830 224.760 144.130 225.760 ;
    END
  END ui_in[1]
  PIN ui_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 140.150 224.760 140.450 225.760 ;
    END
  END ui_in[2]
  PIN ui_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 136.470 224.760 136.770 225.760 ;
    END
  END ui_in[3]
  PIN ui_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 132.790 224.760 133.090 225.760 ;
    END
  END ui_in[4]
  PIN ui_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 129.110 224.760 129.410 225.760 ;
    END
  END ui_in[5]
  PIN ui_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 125.430 224.760 125.730 225.760 ;
    END
  END ui_in[6]
  PIN ui_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 121.750 224.760 122.050 225.760 ;
    END
  END ui_in[7]
  PIN uio_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 118.070 224.760 118.370 225.760 ;
    END
  END uio_in[0]
  PIN uio_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 114.390 224.760 114.690 225.760 ;
    END
  END uio_in[1]
  PIN uio_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 110.710 224.760 111.010 225.760 ;
    END
  END uio_in[2]
  PIN uio_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 107.030 224.760 107.330 225.760 ;
    END
  END uio_in[3]
  PIN uio_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 103.350 224.760 103.650 225.760 ;
    END
  END uio_in[4]
  PIN uio_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 99.670 224.760 99.970 225.760 ;
    END
  END uio_in[5]
  PIN uio_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 95.990 224.760 96.290 225.760 ;
    END
  END uio_in[6]
  PIN uio_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 92.310 224.760 92.610 225.760 ;
    END
  END uio_in[7]
  PIN uio_oe[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 29.750 224.760 30.050 225.760 ;
    END
  END uio_oe[0]
  PIN uio_oe[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 26.070 224.760 26.370 225.760 ;
    END
  END uio_oe[1]
  PIN uio_oe[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 22.390 224.760 22.690 225.760 ;
    END
  END uio_oe[2]
  PIN uio_oe[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 18.710 224.760 19.010 225.760 ;
    END
  END uio_oe[3]
  PIN uio_oe[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 15.030 224.760 15.330 225.760 ;
    END
  END uio_oe[4]
  PIN uio_oe[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 11.350 224.760 11.650 225.760 ;
    END
  END uio_oe[5]
  PIN uio_oe[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 7.670 224.760 7.970 225.760 ;
    END
  END uio_oe[6]
  PIN uio_oe[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 3.990 224.760 4.290 225.760 ;
    END
  END uio_oe[7]
  PIN uio_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 59.190 224.760 59.490 225.760 ;
    END
  END uio_out[0]
  PIN uio_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 55.510 224.760 55.810 225.760 ;
    END
  END uio_out[1]
  PIN uio_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 51.830 224.760 52.130 225.760 ;
    END
  END uio_out[2]
  PIN uio_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 48.150 224.760 48.450 225.760 ;
    END
  END uio_out[3]
  PIN uio_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 44.470 224.760 44.770 225.760 ;
    END
  END uio_out[4]
  PIN uio_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 40.790 224.760 41.090 225.760 ;
    END
  END uio_out[5]
  PIN uio_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 37.110 224.760 37.410 225.760 ;
    END
  END uio_out[6]
  PIN uio_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 33.430 224.760 33.730 225.760 ;
    END
  END uio_out[7]
  PIN uo_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 88.630 224.760 88.930 225.760 ;
    END
  END uo_out[0]
  PIN uo_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 84.950 224.760 85.250 225.760 ;
    END
  END uo_out[1]
  PIN uo_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 81.270 224.760 81.570 225.760 ;
    END
  END uo_out[2]
  PIN uo_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 77.590 224.760 77.890 225.760 ;
    END
  END uo_out[3]
  PIN uo_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 73.910 224.760 74.210 225.760 ;
    END
  END uo_out[4]
  PIN uo_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 70.230 224.760 70.530 225.760 ;
    END
  END uo_out[5]
  PIN uo_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 66.550 224.760 66.850 225.760 ;
    END
  END uo_out[6]
  PIN uo_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 62.870 224.760 63.170 225.760 ;
    END
  END uo_out[7]
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1.000 5.000 2.500 220.760 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 49.000 5.000 50.500 220.760 ;
    END
  END VGND
  OBS
      LAYER nwell ;
        RECT 85.850 83.495 89.560 100.755 ;
        RECT 100.875 96.805 103.650 118.465 ;
        RECT 84.510 80.095 89.560 83.495 ;
        RECT 85.850 43.085 89.560 80.095 ;
        RECT 108.455 63.635 113.020 118.860 ;
        RECT 107.190 60.235 113.020 63.635 ;
        RECT 108.455 18.195 113.020 60.235 ;
      LAYER li1 ;
        RECT 109.640 118.805 111.970 118.975 ;
        RECT 102.300 118.135 102.470 118.155 ;
        RECT 101.205 115.255 102.470 118.135 ;
        RECT 98.730 113.755 102.470 115.255 ;
        RECT 84.905 80.445 85.665 83.135 ;
        RECT 86.245 43.400 86.415 100.440 ;
        RECT 87.035 43.400 87.205 100.440 ;
        RECT 87.825 43.400 87.995 100.440 ;
        RECT 88.435 78.255 89.195 100.385 ;
        RECT 101.205 97.135 102.470 113.755 ;
        RECT 102.300 97.115 102.470 97.135 ;
        RECT 103.090 96.810 103.260 118.155 ;
        RECT 106.300 110.030 107.060 110.615 ;
        RECT 102.950 96.430 103.375 96.810 ;
        RECT 100.945 95.630 101.565 96.180 ;
        RECT 102.300 95.630 102.470 95.650 ;
        RECT 100.935 95.200 102.470 95.630 ;
        RECT 102.300 95.180 102.470 95.200 ;
        RECT 103.090 95.180 103.260 96.430 ;
        RECT 100.130 93.755 100.635 94.255 ;
        RECT 102.510 94.090 103.045 94.550 ;
        RECT 104.225 93.755 105.735 97.250 ;
        RECT 96.230 89.255 97.730 90.755 ;
        RECT 95.250 85.365 95.420 88.805 ;
        RECT 96.040 85.365 96.210 88.805 ;
        RECT 93.710 84.795 94.340 85.265 ;
        RECT 93.920 84.285 94.090 84.795 ;
        RECT 94.805 84.340 95.305 84.755 ;
        RECT 93.400 83.895 94.130 84.285 ;
        RECT 88.435 75.755 92.230 78.255 ;
        RECT 88.435 43.470 89.195 75.755 ;
        RECT 93.400 75.365 93.570 83.895 ;
        RECT 94.190 74.955 94.360 83.405 ;
        RECT 94.980 75.365 95.150 84.340 ;
        RECT 95.805 79.255 96.655 83.315 ;
        RECT 95.805 78.255 98.730 79.255 ;
        RECT 95.805 75.450 96.655 78.255 ;
        RECT 99.900 75.645 100.070 92.685 ;
        RECT 100.690 75.645 100.860 92.685 ;
        RECT 103.290 88.845 103.460 92.885 ;
        RECT 104.080 88.845 104.250 92.885 ;
        RECT 102.730 84.250 104.730 86.255 ;
        RECT 106.190 84.305 106.360 109.345 ;
        RECT 106.980 84.305 107.150 109.345 ;
        RECT 106.230 81.760 107.235 82.755 ;
        RECT 96.145 74.955 96.315 75.450 ;
        RECT 94.190 74.785 96.315 74.955 ;
        RECT 107.585 60.585 108.345 63.275 ;
        RECT 89.230 37.515 90.230 39.255 ;
        RECT 92.340 39.015 94.510 39.365 ;
        RECT 95.010 39.015 97.170 39.365 ;
        RECT 92.340 37.515 94.420 39.015 ;
        RECT 89.230 37.330 94.420 37.515 ;
        RECT 95.110 37.930 97.170 39.015 ;
        RECT 95.110 37.330 97.175 37.930 ;
        RECT 89.230 36.980 94.515 37.330 ;
        RECT 95.015 37.000 97.175 37.330 ;
        RECT 98.230 37.000 99.230 39.255 ;
        RECT 95.015 36.980 99.235 37.000 ;
        RECT 89.230 36.430 94.420 36.980 ;
        RECT 92.340 35.225 94.420 36.430 ;
        RECT 95.110 36.150 99.235 36.980 ;
        RECT 95.110 35.780 97.175 36.150 ;
        RECT 95.110 35.225 97.170 35.780 ;
        RECT 92.340 34.875 94.500 35.225 ;
        RECT 95.000 34.875 97.170 35.225 ;
        RECT 89.550 32.450 90.625 33.300 ;
        RECT 92.340 32.975 94.420 34.875 ;
        RECT 95.110 32.975 97.170 34.875 ;
        RECT 92.340 32.625 94.500 32.975 ;
        RECT 95.000 32.625 97.170 32.975 ;
        RECT 92.340 30.430 94.005 32.625 ;
        RECT 95.110 32.615 97.170 32.625 ;
        RECT 108.850 18.505 109.020 118.545 ;
        RECT 109.640 18.205 109.810 118.805 ;
        RECT 110.430 18.505 110.600 118.545 ;
        RECT 111.800 118.440 111.970 118.805 ;
        RECT 110.945 77.245 112.690 118.440 ;
        RECT 110.945 75.755 115.240 77.245 ;
        RECT 110.945 27.755 112.690 75.755 ;
        RECT 110.945 26.255 115.230 27.755 ;
        RECT 110.945 18.850 112.690 26.255 ;
        RECT 111.720 18.205 111.890 18.850 ;
        RECT 109.640 18.035 111.890 18.205 ;
      LAYER mcon ;
        RECT 99.015 114.025 99.965 114.990 ;
        RECT 85.100 81.325 85.450 81.765 ;
        RECT 86.245 43.480 86.415 100.360 ;
        RECT 87.035 43.480 87.205 100.360 ;
        RECT 87.825 43.480 87.995 100.360 ;
        RECT 102.300 97.195 102.470 118.075 ;
        RECT 103.090 97.195 103.260 118.075 ;
        RECT 106.440 110.180 106.935 110.545 ;
        RECT 101.015 95.720 101.360 96.050 ;
        RECT 102.300 95.260 102.470 95.570 ;
        RECT 103.090 95.260 103.260 95.570 ;
        RECT 104.690 95.235 105.275 95.790 ;
        RECT 100.210 93.855 100.555 94.175 ;
        RECT 102.590 94.170 102.965 94.470 ;
        RECT 96.480 89.520 97.485 90.540 ;
        RECT 95.250 85.445 95.420 88.725 ;
        RECT 96.040 85.445 96.210 88.725 ;
        RECT 93.850 84.875 94.230 85.175 ;
        RECT 94.870 84.400 95.250 84.670 ;
        RECT 93.400 75.445 93.570 83.325 ;
        RECT 94.190 75.445 94.360 83.325 ;
        RECT 94.980 75.445 95.150 83.325 ;
        RECT 97.970 78.430 98.545 79.060 ;
        RECT 99.900 75.725 100.070 92.605 ;
        RECT 100.690 75.725 100.860 92.605 ;
        RECT 103.290 88.925 103.460 92.805 ;
        RECT 104.080 88.925 104.250 92.805 ;
        RECT 103.325 85.475 104.070 86.070 ;
        RECT 106.190 84.385 106.360 109.265 ;
        RECT 106.980 84.385 107.150 109.265 ;
        RECT 106.465 82.005 107.035 82.555 ;
        RECT 107.780 61.465 108.130 61.905 ;
        RECT 98.455 38.505 99.025 39.075 ;
        RECT 89.650 32.545 90.500 33.200 ;
        RECT 92.615 30.600 93.680 31.265 ;
        RECT 108.850 18.585 109.020 118.465 ;
        RECT 109.640 18.585 109.810 118.465 ;
        RECT 110.430 18.585 110.600 118.465 ;
        RECT 114.065 76.170 114.910 76.960 ;
        RECT 114.045 26.520 114.900 27.420 ;
      LAYER met1 ;
        RECT 106.350 119.350 111.230 119.950 ;
        RECT 98.730 113.755 100.230 115.255 ;
        RECT 86.215 102.575 95.235 102.935 ;
        RECT 86.215 100.420 86.450 102.575 ;
        RECT 87.795 102.045 94.210 102.405 ;
        RECT 85.020 81.255 85.540 81.875 ;
        RECT 86.215 43.420 86.445 100.420 ;
        RECT 86.700 42.755 87.535 100.550 ;
        RECT 87.795 43.420 88.025 102.045 ;
        RECT 93.850 85.265 94.210 102.045 ;
        RECT 94.875 94.255 95.235 102.575 ;
        RECT 102.270 97.135 102.500 118.135 ;
        RECT 103.060 97.135 103.290 118.135 ;
        RECT 106.350 110.615 106.950 119.350 ;
        RECT 110.630 118.525 111.230 119.350 ;
        RECT 106.300 110.030 107.060 110.615 ;
        RECT 100.945 95.630 101.440 96.180 ;
        RECT 102.270 95.200 102.500 95.630 ;
        RECT 103.060 95.200 103.290 95.630 ;
        RECT 94.875 93.755 100.630 94.255 ;
        RECT 102.510 94.090 103.045 94.550 ;
        RECT 104.225 93.755 105.735 97.250 ;
        RECT 94.875 88.785 95.235 93.755 ;
        RECT 106.160 92.865 106.390 109.325 ;
        RECT 96.230 89.255 97.730 90.755 ;
        RECT 94.875 85.385 95.450 88.785 ;
        RECT 96.010 87.255 96.240 88.785 ;
        RECT 96.010 86.255 98.230 87.255 ;
        RECT 96.010 85.385 96.240 86.255 ;
        RECT 93.710 84.795 94.340 85.265 ;
        RECT 94.875 84.755 95.235 85.385 ;
        RECT 94.805 84.340 95.305 84.755 ;
        RECT 90.090 75.755 92.230 78.255 ;
        RECT 93.370 75.385 93.600 83.385 ;
        RECT 94.160 75.385 94.390 83.385 ;
        RECT 94.950 75.385 95.180 83.385 ;
        RECT 99.230 79.255 100.100 92.665 ;
        RECT 97.730 78.255 100.100 79.255 ;
        RECT 99.230 75.665 100.100 78.255 ;
        RECT 100.660 82.755 101.730 92.665 ;
        RECT 102.730 88.865 103.490 92.865 ;
        RECT 104.050 91.255 106.390 92.865 ;
        RECT 104.050 90.755 104.310 91.255 ;
        RECT 106.130 90.755 106.390 91.255 ;
        RECT 104.050 90.255 106.390 90.755 ;
        RECT 104.050 89.755 104.310 90.255 ;
        RECT 106.130 89.755 106.390 90.255 ;
        RECT 104.050 88.865 106.390 89.755 ;
        RECT 102.730 87.755 103.260 88.865 ;
        RECT 102.730 84.250 104.730 87.755 ;
        RECT 106.160 84.325 106.390 88.865 ;
        RECT 106.950 107.755 107.180 109.325 ;
        RECT 106.950 106.255 107.970 107.755 ;
        RECT 106.950 90.755 107.180 106.255 ;
        RECT 106.950 89.255 108.030 90.755 ;
        RECT 106.950 84.325 107.180 89.255 ;
        RECT 100.660 81.760 107.235 82.755 ;
        RECT 100.660 75.665 101.730 81.760 ;
        RECT 100.890 74.255 101.730 75.665 ;
        RECT 107.700 61.395 108.220 62.015 ;
        RECT 108.820 47.390 109.050 118.525 ;
        RECT 106.220 42.755 109.050 47.390 ;
        RECT 86.700 40.685 109.050 42.755 ;
        RECT 98.230 38.255 99.230 39.255 ;
        RECT 106.220 35.250 109.050 40.685 ;
        RECT 89.550 32.450 90.625 33.300 ;
        RECT 92.340 30.430 94.005 31.490 ;
        RECT 108.820 18.525 109.050 35.250 ;
        RECT 109.610 18.525 109.840 118.525 ;
        RECT 110.400 18.525 111.230 118.525 ;
        RECT 113.730 75.755 115.240 77.245 ;
        RECT 113.730 26.255 115.230 27.755 ;
      LAYER via ;
        RECT 99.015 114.025 99.965 114.990 ;
        RECT 85.100 81.325 85.450 81.765 ;
        RECT 101.015 95.720 101.360 96.050 ;
        RECT 104.690 95.235 105.275 95.790 ;
        RECT 102.590 94.170 102.965 94.470 ;
        RECT 96.480 89.520 97.485 90.540 ;
        RECT 97.425 86.460 98.040 87.060 ;
        RECT 90.525 76.100 91.880 77.850 ;
        RECT 97.970 78.430 98.545 79.060 ;
        RECT 104.690 91.615 105.590 92.565 ;
        RECT 103.515 86.500 104.440 87.510 ;
        RECT 107.330 106.595 107.820 107.535 ;
        RECT 107.330 89.350 107.860 90.565 ;
        RECT 101.040 74.370 101.600 74.930 ;
        RECT 107.780 61.465 108.130 61.905 ;
        RECT 98.455 38.505 99.025 39.075 ;
        RECT 89.650 32.545 90.500 33.200 ;
        RECT 92.615 30.600 93.680 31.265 ;
        RECT 114.065 76.170 114.910 76.960 ;
        RECT 114.045 26.520 114.900 27.420 ;
      LAYER met2 ;
        RECT 79.840 115.255 81.825 120.040 ;
        RECT 79.840 113.755 100.230 115.255 ;
        RECT 79.840 107.755 81.825 113.755 ;
        RECT 79.840 106.255 107.970 107.755 ;
        RECT 79.840 90.755 81.825 106.255 ;
        RECT 104.225 96.180 105.735 97.250 ;
        RECT 117.725 96.180 119.710 119.970 ;
        RECT 100.945 95.760 119.710 96.180 ;
        RECT 100.945 95.630 101.565 95.760 ;
        RECT 91.060 92.450 91.895 92.755 ;
        RECT 102.510 92.450 103.045 94.550 ;
        RECT 104.225 93.755 105.735 95.760 ;
        RECT 91.060 91.915 103.045 92.450 ;
        RECT 91.060 91.725 91.895 91.915 ;
        RECT 104.395 91.310 106.005 92.820 ;
        RECT 79.840 89.255 108.030 90.755 ;
        RECT 79.840 82.315 81.825 89.255 ;
        RECT 117.725 87.755 119.710 95.760 ;
        RECT 97.230 86.255 98.230 87.255 ;
        RECT 103.260 86.255 119.710 87.755 ;
        RECT 79.840 80.805 85.640 82.315 ;
        RECT 79.840 78.255 81.825 80.805 ;
        RECT 117.725 79.255 119.710 86.255 ;
        RECT 97.730 78.255 119.710 79.255 ;
        RECT 79.840 77.245 92.230 78.255 ;
        RECT 79.840 75.755 115.240 77.245 ;
        RECT 79.840 62.455 81.825 75.755 ;
        RECT 100.890 74.255 101.730 75.020 ;
        RECT 79.840 60.945 108.320 62.455 ;
        RECT 79.840 27.755 81.825 60.945 ;
        RECT 98.230 38.255 99.230 39.255 ;
        RECT 89.550 32.450 90.625 33.300 ;
        RECT 92.340 30.430 94.005 31.490 ;
        RECT 79.840 26.255 115.230 27.755 ;
        RECT 79.840 18.100 81.825 26.255 ;
        RECT 117.725 18.030 119.710 78.255 ;
      LAYER via2 ;
        RECT 91.250 91.925 91.710 92.575 ;
        RECT 104.690 91.615 105.590 92.565 ;
        RECT 97.425 86.460 98.040 87.060 ;
        RECT 101.040 74.370 101.600 74.930 ;
        RECT 98.455 38.505 99.025 39.075 ;
        RECT 89.650 32.545 90.500 33.200 ;
        RECT 92.615 30.600 93.680 31.265 ;
        RECT 80.130 18.465 81.515 19.795 ;
        RECT 118.290 18.360 119.140 19.190 ;
      LAYER met3 ;
        RECT 86.570 94.655 113.630 125.055 ;
        RECT 91.060 92.570 91.895 92.755 ;
        RECT 86.295 91.920 91.895 92.570 ;
        RECT 86.295 25.775 86.945 91.920 ;
        RECT 91.060 91.725 91.895 91.920 ;
        RECT 104.395 92.690 113.630 94.655 ;
        RECT 104.395 91.690 115.120 92.690 ;
        RECT 104.395 91.310 106.005 91.690 ;
        RECT 97.230 73.730 98.230 87.255 ;
        RECT 100.890 74.255 101.730 75.020 ;
        RECT 91.295 43.330 105.155 73.730 ;
        RECT 114.120 39.255 115.120 91.690 ;
        RECT 98.230 38.255 115.120 39.255 ;
        RECT 89.550 32.450 90.625 33.300 ;
        RECT 92.340 30.430 94.005 31.490 ;
        RECT 86.000 22.255 87.245 25.775 ;
        RECT 79.835 18.095 81.830 20.115 ;
        RECT 117.720 18.030 119.720 19.320 ;
      LAYER via3 ;
        RECT 113.210 94.795 113.530 124.915 ;
        RECT 101.040 74.370 101.600 74.930 ;
        RECT 104.735 43.470 105.055 73.590 ;
        RECT 103.200 38.435 103.940 39.135 ;
        RECT 89.650 32.545 90.500 33.200 ;
        RECT 92.615 30.600 93.680 31.265 ;
        RECT 86.120 22.500 87.090 23.360 ;
        RECT 80.130 18.465 81.515 19.795 ;
        RECT 118.290 18.360 119.140 19.190 ;
      LAYER met4 ;
        RECT 86.965 111.415 111.775 124.660 ;
        RECT 82.625 109.400 111.775 111.415 ;
        RECT 82.625 34.810 84.640 109.400 ;
        RECT 86.965 95.050 111.775 109.400 ;
        RECT 113.130 94.715 113.610 124.995 ;
        RECT 100.890 73.335 101.730 75.020 ;
        RECT 91.690 43.725 103.300 73.335 ;
        RECT 104.655 43.390 105.135 73.670 ;
        RECT 76.845 34.015 84.640 34.810 ;
        RECT 48.175 30.110 49.000 34.015 ;
        RECT 50.500 30.110 84.640 34.015 ;
        RECT 76.845 30.105 82.975 30.110 ;
        RECT 89.550 29.245 90.625 33.300 ;
        RECT 92.340 30.430 97.150 31.450 ;
        RECT 89.550 28.105 92.745 29.245 ;
        RECT 85.925 20.340 87.380 23.630 ;
        RECT 59.885 18.090 81.925 20.110 ;
        RECT 60.390 2.175 61.405 18.090 ;
        RECT 86.110 6.740 87.190 20.340 ;
        RECT 91.310 15.605 92.730 28.105 ;
        RECT 90.090 14.540 92.730 15.605 ;
        RECT 68.000 5.660 87.190 6.740 ;
        RECT 46.160 1.575 61.405 2.175 ;
        RECT 46.160 1.000 46.760 1.575 ;
        RECT 60.390 1.370 61.405 1.575 ;
        RECT 68.240 1.000 68.840 5.660 ;
        RECT 90.320 1.000 90.920 14.540 ;
        RECT 91.310 14.360 92.730 14.540 ;
        RECT 95.845 9.650 97.145 30.430 ;
        RECT 102.995 13.950 104.110 39.385 ;
        RECT 117.720 19.310 119.710 19.320 ;
        RECT 117.720 18.090 157.470 19.310 ;
        RECT 117.720 18.030 119.710 18.090 ;
        RECT 102.995 12.835 135.340 13.950 ;
        RECT 95.845 8.580 113.235 9.650 ;
        RECT 95.845 8.465 97.145 8.580 ;
        RECT 112.400 1.000 113.000 8.580 ;
        RECT 134.480 1.000 135.080 12.835 ;
        RECT 156.560 1.000 157.160 18.090 ;
  END
END tt_um_duk_opamp
END LIBRARY

